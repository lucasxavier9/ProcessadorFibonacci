module adder (
    input logic [7:0] a, b,
    output logic [7:0] s
);
   assign s = a + b;
   
endmodule